module adder(input a,b,output c);

    assign c==a+b;

endmodule
